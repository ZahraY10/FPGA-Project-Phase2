library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.math_real.all;
use IEEE.numeric_std.all;

library work;
use work.neurals_utils.all;

entity input is
    Port (
        xt: in matrix_1_4;
        ht_1: in matrix_1_8;
        i: out matrix_1_8
    );
end input;

architecture Behavioral of input is

    signal wi: matrix_4_8 := (
    (0.13965783,-0.04775485,0.34143683,0.28217432,0.05485592,0.5929077,-0.14488743,0.0269083),
    (-0.26471546,0.21732531,-0.63501525,-0.5341712,0.4722219,0.1886938,0.16185956,-0.1487629),
    (0.3210674,0.32791585,0.24699497,-0.19182979,0.21832567,0.22613047,0.1668725,-0.10851475), 
    (0.09162864,-0.22094683,-0.7704977,-0.27422312,-0.5308995,-0.19721255,-0.10660882,-0.28635386));

    signal ui: matrix_8_8 := (
    (-0.22540611,-0.07725633,-0.04325512,-0.04499104,-0.32806206,-0.04144218,-0.03638914,0.03160138),
    (0.18012986,-0.29333568,0.00671834,-0.16674466,-0.34768414,0.01304776,-0.06656786,-0.33698344),
    (0.35989136,-0.16509496,-0.07809209,-0.02823459,-0.6466683,0.03439626,-0.02917804,0.06093279),
    (0.20940925,0.38939223,0.02142915,0.06047469,0.19592714,0.50517815,0.14237255,0.48360968),
    (0.02413642,0.16279134,0.02921131,0.4190974,-0.31731865,-0.16067709,0.34781075,0.07166091),
    (-0.07821875,0.14518033,-0.35107407,-0.02979031,0.25414816,-0.37739775,0.45078024,0.20540176),
    (0.11960886,-0.00708573,-0.01591504,-0.0124966,0.23815277,0.15988702,-0.10813737,0.17890273),
    (0.28208584,0.28524047,-0.11078832,0.05000078,0.62929094,0.03044126,0.37248662,0.19190663));
    
    signal bi: matrix_1_8 := (
      0.22003067,
      0.3905463,
      0.21280797,
      0.22266074,
      0.5750835,
      0.5361282,
      0.19412729,
      0.18189429);
    
    signal xt_wi: matrix_1_8 := (others => 0.0);
    signal ht_1_ui: matrix_1_8 := (others => 0.0);
         
     
begin

    process
    variable temp : real := 0.0;
    begin
        F1: for t in 0 to 7 loop
            F2: for j in 0 to 3 loop
                temp := xt(j) * wi(j, t);
                xt_wi(t) <= xt_wi(t) + temp;  
            end loop F2;
        end loop F1;
        
        F3: for t in 0 to 7 loop
            F4: for j in 0 to 7 loop
                temp := ht_1(j) * ui(j, t);
                ht_1_ui(t) <= ht_1_ui(t) + temp;  
            end loop F4;
        end loop F3;
        
        F5: for t in 0 to 7 loop
            temp := bi(t) + ht_1_ui(t);
            i(t) <= temp + xt_wi(t);
        end loop F5;
            
    end process;
end Behavioral;
