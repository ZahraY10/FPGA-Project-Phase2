library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.math_real.all;
use IEEE.numeric_std.all;

library work;
use work.neurals_utils.all;

entity output is
    Port (
        xt: in matrix_1_4;
        ht_1: in matrix_1_8;
        o: out matrix_1_8
    );
end output;

architecture Behavioral of output is

    signal wo: matrix_4_8 := (
    (0.81262547,0.3234628,0.7666596,-0.14796887,1.0295157,0.5463878,-0.2399153,-0.29666474),
    (0.7540123,-0.07887857,-0.72580874,-0.41807404,0.07835332,-0.90355235,-0.07551592,-0.37188026),
    (0.46900183,0.04062076,1.0506912,-0.20407581,0.53115785,0.49669996,0.15442692,0.02013548), 
    (-0.32798606,0.03164255,-0.6752109,-0.5345587,-0.82918984,0.0482377,0.05022579,0.12873164));

    signal uo: matrix_8_8 := (
    (-0.1564388,0.060792,-0.25346947,-0.21916276,-0.05961246,0.16500823,0.07056013,-0.04299608),
    (-0.10268968,-0.16318482,-0.0763059,-0.14473884,-0.32715902,-0.3284195,0.01457982,-0.21989729),
    (0.4014409,-0.20964584,0.12663233,0.15928917,0.06926352,0.0872872,0.09628288,0.20289727),
    (0.31969658,0.48952508,-0.06890938,0.04971746,0.4850268,0.77359366,0.04772833,0.00763122),
    (-0.21406649,0.3851055,0.06895181,-0.09096608,0.2268963,0.02800295,-0.26645523,0.09101521),
    (-0.23577942,0.40463912,-0.02379321,0.12271876,0.20454015,0.3340834,0.20872128,0.23313737),
    (0.36070636,-0.08882497,0.1167473,-0.09869172,0.3148002,0.41594255,-0.1424936,-0.13277136),
    (-0.09099162,-0.14975166,0.14469796,-0.09419464,0.34336716,0.45454732,-0.19643505,0.19911067));
    
    signal bo: matrix_1_8 := (
      0.215092,
      0.48508435,
      0.2803704,
      0.26674628,
      0.60106176,
      0.65973246,
      0.22069259,
      0.21072803);
    
    signal xt_wo: matrix_1_8 := (others => 0.0);
    signal ht_1_uo: matrix_1_8 := (others => 0.0);
         
     
begin

    process
    variable temp : real := 0.0;
    begin
        F1: for i in 0 to 7 loop
            F2: for j in 0 to 3 loop
                temp := xt(j) * wo(j, i);
                xt_wo(i) <= xt_wo(i) + temp;  
            end loop F2;
        end loop F1;
        
        F3: for i in 0 to 7 loop
            F4: for j in 0 to 7 loop
                temp := ht_1(j) * uo(j, i);
                ht_1_uo(i) <= ht_1_uo(i) + temp;  
            end loop F4;
        end loop F3;
        
        F5: for i in 0 to 7 loop
            temp := bo(i) + ht_1_uo(i);
            o(i) <= temp + xt_wo(i);
        end loop F5;
            
    end process;
end Behavioral;
