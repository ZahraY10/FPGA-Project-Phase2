library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.math_real.all;
use IEEE.numeric_std.all;

library work;
use work.neurals_utils.all;

entity candidate is
    Port (
        xt: in matrix_1_4;
        ht_1: in matrix_1_8;
        cnd: out matrix_1_8
    );
end candidate;

architecture Behavioral of candidate is

    signal wc: matrix_4_8 := (
    (-0.21440436,0.58637863,-0.07314462,0.6577152,-0.8901406,-0.49870068,0.7506063,-0.14046632),
    (0.08641554,-0.01217922,0.13672125,-0.75612044,0.6853312,-0.2585029,-0.7974984,0.16907303),
    (-0.73499763,0.5950351,-0.20747943,0.3708285,-0.76652896,-0.57712734,0.54822814,-0.24967012), 
    (0.25779077,-0.60224974,-0.2717871,-0.18705575,0.82094723,0.6652274,-0.21723086,0.17782894));

    signal uc: matrix_8_8 := (
    (0.24807113,-0.18499182,-0.48871857,-0.05675852,0.1581574,0.4236816,-0.22095923,0.12871744),
    (-0.177079,0.4365895,-0.10886224,-0.2711792,0.06320903,-0.3596882,0.03018917,-0.16216652),
    (-0.01938948,0.1877461,0.21442765,-0.18974146,-0.19947451,-0.09283099,-0.42934605,-0.09511761),
    (-0.52744734,0.32326484,0.28837425,0.3303778,-0.264037,-0.11096267,0.25911146,-0.30506),
    (0.22532704,-0.1567047,-0.33357525,-0.03777692,-0.03376415,0.5673492,0.03478994,0.02179503),
    (-0.2492082,-0.15948121,-0.26482478,-0.03805209,-0.00448201,0.07136463,-0.11671741,0.22851901),
    (-0.12679164,0.5482961,-0.05207148,0.03086551,-0.4302712,-0.49658602,0.06617329,-0.5270848),
    (0.21930438,-0.07057948,-0.04036796,-0.1382596,-0.00983683,0.09509208,0.2272774,0.22204381));
    
    signal bc: matrix_1_8 := (
     -0.05570378,
     -0.00401851,
     0.1789396,
     -0.00899142,
     -0.02097004,
     -0.00503316,
     0.02325593,
     0.00892116);
    
    signal xt_wc: matrix_1_8 := (others => 0.0);
    signal ht_1_uc: matrix_1_8 := (others => 0.0);
         
     
begin

    process
    variable temp : real := 0.0;
    begin
        F1: for i in 0 to 7 loop
            F2: for j in 0 to 3 loop
                temp := xt(j) * wc(j, i);
                xt_wc(i) <= xt_wc(i) + temp;  
            end loop F2;
        end loop F1;
        
        F3: for i in 0 to 7 loop
            F4: for j in 0 to 7 loop
                temp := ht_1(j) * uc(j, i);
                ht_1_uc(i) <= ht_1_uc(i) + temp;  
            end loop F4;
        end loop F3;
        
        F5: for i in 0 to 7 loop
            temp := bc(i) + ht_1_uc(i);
            cnd(i) <= temp + xt_wc(i);
        end loop F5;
            
    end process;
end Behavioral;
